/////////////////////////////////////////PC_MODULE///////////////////////////////////////////////////////////////
module PC
(
    input clk,res,
    input [31:0] in,
    output reg [31:0] out
);
 
  always@(posedge clk or posedge res) begin
    if(res)
      out<=32'b0;
    else
      out<=in;
  end

endmodule
//////////////////////////////////////////////////////////////////////////////////////////////////////////////
